`timescale 1ns / 1ps
`default_nettype none

module intersection_detector(
    input wire clk_pixel_in,
    input wire rst_in,
    input wire is_attacking,
    input wire [10:0] saber_start_x,
    input wire [9:0] saber_start_y,
    input wire [10:0] saber_current_x,
    input wire [9:0] saber_current_y,
    input location_t opponent,
    output logic is_intersecting
  );

  
  
endmodule

`default_nettype wire
